module AlteraProject(A, B, C);

output A;
input B, C;

assign A = B | C;

endmodule

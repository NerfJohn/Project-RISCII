/*
 * ImmBlock.v
 *
 * "Generates immediate value based on given opcode"
 */
module ImmBlock (
	// Input instruction connection.
	input  [7:0]  i_instrImm,
	input  [3:0]  i_instrOpcode,
	
	// Output immediate connection.
	output [15:0] o_genImm
);

/*
 * TODO- desc.
 */

////////////////////////////////////////////////////////////////////////////////
// -- Internal Signals/Wires -- //
////////////////////////////////////////////////////////////////////////////////

// Computed controls based on opcode.
wire        isSize8;
wire        doShift;

// Base selection wires.
wire [15:0] baseImm;

// Length resolution wires.
wire [15:0] immSized;
	
////////////////////////////////////////////////////////////////////////////////
// -- Connections/Comb Logic -- //
////////////////////////////////////////////////////////////////////////////////

//------------------------------------------------------------------------------
// Compute opcode based controls.
//assign isSize6 = ~i_instrOpcode[3] & ~i_instrOpcode[1];
assign isSize8 = ~i_instrOpcode[2] &  i_instrOpcode[1] & ~i_instrOpcode[0];
assign doShift = ~i_instrOpcode[3];

//------------------------------------------------------------------------------
// Compute base immediate.
Mux2 M0[15:0] (
	.A({{8{i_instrImm[7]}}, i_instrImm}),       // 8-bit imm? generate int8
	.B({{11{i_instrImm[4]}}, i_instrImm[4:0]}), // No?        generate int5
	.S(isSize8),
	.Y(baseImm)
);

//------------------------------------------------------------------------------
// Drive generated immediate (shifting for control opcodes).
Mux2 M1[15:0] (
	.A({baseImm[14:0], 1'b0}), // Shift? return base left shifted by 1 bit
	.B(baseImm),               // No?    return base
	.S(doShift),
	.Y(o_genImm)
);

endmodule

module timer_16b(busAddr, busData, busEn, busWr,	// Bus Access
                 sigIntr, clk2,							// Special Signals
					  clk, rstn,								// Common Signals
					  TEST_cnt, TEST_ctrl					// Test points (TODO- Remove)
);
					  
/* TODO- Module Desc. */

// -- Signals -- //

// Common CLK/RST lines.
input clk, rstn;

// Special signals.
input clk2;				// 2nd selectable clock source for timer
output sigIntr;		// Interrupt signal generated by overflow

// Bus signals.
input[1:0] busAddr;	// Sub-address of timer's internal registers
input busEn;			// Enable to trigger read/write
input busWr;			// Signal to distinguish read/write requests
inout[15:0] busData;	// Data used to write in/read out data

// TEST signals: TODO- remove.
output[15:0] TEST_cnt, TEST_ctrl;

// Basic loop of timer.
wire[15:0] incIn, incOut, valIn;

// -- Instances -- //

// Internal Registers- value, control, and max register.
dff_en iVR[15:0] (.D(valIn), .Q(incIn), .en(~busEn | busWr), .clk(clk), .rstn(rstn));

// Adder for actual incrementing.
add_16b iINC (.src1(incIn), .src2(16'b0), .cin(1'b1), .sum(incOut), .cout(/*NC*/));

// Write selection- allow bus to write to value register.
mux2 iMUX0[15:0] (.A(busData), .B(incOut), .sel(busEn), .out(valIn));

// -- Raw Logic -- //

// Tristate input to bus.
assign busData = (busEn & ~busWr) ? incIn : 16'bz;

// TEST signals: TODO- remove.
assign TEST_cnt = incIn;

// (TODO- implement.)
assign sigIntr = 0;
assign TEST_ctrl = 0;

/*
// Intermediate signals.
wire selClk;
wire[7:0] crOut;
wire[15:0] vrOut, mrOut;
wire[15:0] vrIn;
wire[3:0] psIn, psOut;

// -- Instances -- //

// Internal Registers- value, control, and max register.
mux2 iMUX0[15:0] (.A(busData), .B(), .sel(busEn), .out(vrIn));
dff_en iVR[15:0] (.D(vrIn), .Q(vrOut), .en(), .clk(selClk), .rstn(rstn));
dff_en iCR[7:0]  (.D(), .Q(crOut), .en(), .clk(selClk), .rstn(rstn));
dff_en iMR[15:0] (.D(), .Q(mrOut), .en(), .clk(selClk), .rstn(rstn));

// Prescale "counter" register- resets on prescale and control register write.
mux2 iMUX1[3:0] (.A(), .B(), .sel(), .out(psIn));
myDff iPSR[3:0] (.D(psIn), .Q(psOut), .clk(selClk), .rstn(rstn));

// Adders- one for prescaling, the other for actual incrementing.
add_1b iPSA[3:0] (.A(), .B(), .Cin(), .S(), .Cout());
add_16b iINC (.src1(), .src2(), .cin(), .sum(), .cout());

// Clock selection- runs internal registers when bus overrides for read/write.
mux2 iMUX2 (.A(clk2), .B(clk), .sel(crOut[1] & ~busEn), .out(selClk));

// -- Raw Logic -- //
*/

endmodule

library verilog;
use verilog.vl_types.all;
entity sampleCode is
end sampleCode;
